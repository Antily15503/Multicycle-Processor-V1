module cpu 

sudo apt install cpu

endmodule